VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_user_project
  CLASS BLOCK ;
  FOREIGN tiny_user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 14.320 150.000 14.920 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 95.920 150.000 96.520 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 104.080 150.000 104.680 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 112.240 150.000 112.840 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 120.400 150.000 121.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 128.560 150.000 129.160 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 146.000 146.650 150.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 146.000 130.090 150.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 146.000 113.530 150.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 146.000 96.970 150.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 146.000 80.410 150.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 22.480 150.000 23.080 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 146.000 63.850 150.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 146.000 47.290 150.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 146.000 30.730 150.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 146.000 14.170 150.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 30.640 150.000 31.240 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 38.800 150.000 39.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 46.960 150.000 47.560 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 55.120 150.000 55.720 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 63.280 150.000 63.880 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 71.440 150.000 72.040 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 79.600 150.000 80.200 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 87.760 150.000 88.360 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 19.760 150.000 20.360 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 101.360 150.000 101.960 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 109.520 150.000 110.120 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 117.680 150.000 118.280 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 125.840 150.000 126.440 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 134.000 150.000 134.600 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 146.000 135.610 150.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 146.000 119.050 150.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 146.000 102.490 150.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 146.000 85.930 150.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 146.000 69.370 150.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 27.920 150.000 28.520 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 146.000 52.810 150.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 146.000 36.250 150.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 146.000 19.690 150.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 146.000 3.130 150.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 36.080 150.000 36.680 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 44.240 150.000 44.840 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 52.400 150.000 53.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 60.560 150.000 61.160 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 68.720 150.000 69.320 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 76.880 150.000 77.480 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 85.040 150.000 85.640 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 93.200 150.000 93.800 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 17.040 150.000 17.640 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 98.640 150.000 99.240 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 106.800 150.000 107.400 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 114.960 150.000 115.560 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 123.120 150.000 123.720 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 131.280 150.000 131.880 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 146.000 141.130 150.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 146.000 124.570 150.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 146.000 108.010 150.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 146.000 91.450 150.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 146.000 74.890 150.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 25.200 150.000 25.800 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 146.000 58.330 150.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 146.000 41.770 150.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 146.000 25.210 150.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 146.000 8.650 150.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 33.360 150.000 33.960 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 41.520 150.000 42.120 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 49.680 150.000 50.280 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 57.840 150.000 58.440 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 66.000 150.000 66.600 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.160 150.000 74.760 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 82.320 150.000 82.920 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 90.480 150.000 91.080 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.085 10.640 23.685 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.815 10.640 58.415 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.545 10.640 93.145 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.275 10.640 127.875 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.450 10.640 41.050 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.180 10.640 75.780 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.910 10.640 110.510 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.640 10.640 145.240 138.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 4.210 10.640 145.240 138.960 ;
      LAYER met2 ;
        RECT 3.410 145.720 8.090 146.610 ;
        RECT 8.930 145.720 13.610 146.610 ;
        RECT 14.450 145.720 19.130 146.610 ;
        RECT 19.970 145.720 24.650 146.610 ;
        RECT 25.490 145.720 30.170 146.610 ;
        RECT 31.010 145.720 35.690 146.610 ;
        RECT 36.530 145.720 41.210 146.610 ;
        RECT 42.050 145.720 46.730 146.610 ;
        RECT 47.570 145.720 52.250 146.610 ;
        RECT 53.090 145.720 57.770 146.610 ;
        RECT 58.610 145.720 63.290 146.610 ;
        RECT 64.130 145.720 68.810 146.610 ;
        RECT 69.650 145.720 74.330 146.610 ;
        RECT 75.170 145.720 79.850 146.610 ;
        RECT 80.690 145.720 85.370 146.610 ;
        RECT 86.210 145.720 90.890 146.610 ;
        RECT 91.730 145.720 96.410 146.610 ;
        RECT 97.250 145.720 101.930 146.610 ;
        RECT 102.770 145.720 107.450 146.610 ;
        RECT 108.290 145.720 112.970 146.610 ;
        RECT 113.810 145.720 118.490 146.610 ;
        RECT 119.330 145.720 124.010 146.610 ;
        RECT 124.850 145.720 129.530 146.610 ;
        RECT 130.370 145.720 135.050 146.610 ;
        RECT 135.890 145.720 140.570 146.610 ;
        RECT 141.410 145.720 145.210 146.610 ;
        RECT 3.130 4.915 145.210 145.720 ;
      LAYER met3 ;
        RECT 4.400 140.400 146.000 141.265 ;
        RECT 4.000 138.400 146.000 140.400 ;
        RECT 4.400 137.000 146.000 138.400 ;
        RECT 4.000 135.000 146.000 137.000 ;
        RECT 4.400 133.600 145.600 135.000 ;
        RECT 4.000 132.280 146.000 133.600 ;
        RECT 4.000 131.600 145.600 132.280 ;
        RECT 4.400 130.880 145.600 131.600 ;
        RECT 4.400 130.200 146.000 130.880 ;
        RECT 4.000 129.560 146.000 130.200 ;
        RECT 4.000 128.200 145.600 129.560 ;
        RECT 4.400 128.160 145.600 128.200 ;
        RECT 4.400 126.840 146.000 128.160 ;
        RECT 4.400 126.800 145.600 126.840 ;
        RECT 4.000 125.440 145.600 126.800 ;
        RECT 4.000 124.800 146.000 125.440 ;
        RECT 4.400 124.120 146.000 124.800 ;
        RECT 4.400 123.400 145.600 124.120 ;
        RECT 4.000 122.720 145.600 123.400 ;
        RECT 4.000 121.400 146.000 122.720 ;
        RECT 4.400 120.000 145.600 121.400 ;
        RECT 4.000 118.680 146.000 120.000 ;
        RECT 4.000 118.000 145.600 118.680 ;
        RECT 4.400 117.280 145.600 118.000 ;
        RECT 4.400 116.600 146.000 117.280 ;
        RECT 4.000 115.960 146.000 116.600 ;
        RECT 4.000 114.600 145.600 115.960 ;
        RECT 4.400 114.560 145.600 114.600 ;
        RECT 4.400 113.240 146.000 114.560 ;
        RECT 4.400 113.200 145.600 113.240 ;
        RECT 4.000 111.840 145.600 113.200 ;
        RECT 4.000 111.200 146.000 111.840 ;
        RECT 4.400 110.520 146.000 111.200 ;
        RECT 4.400 109.800 145.600 110.520 ;
        RECT 4.000 109.120 145.600 109.800 ;
        RECT 4.000 107.800 146.000 109.120 ;
        RECT 4.400 106.400 145.600 107.800 ;
        RECT 4.000 105.080 146.000 106.400 ;
        RECT 4.000 104.400 145.600 105.080 ;
        RECT 4.400 103.680 145.600 104.400 ;
        RECT 4.400 103.000 146.000 103.680 ;
        RECT 4.000 102.360 146.000 103.000 ;
        RECT 4.000 101.000 145.600 102.360 ;
        RECT 4.400 100.960 145.600 101.000 ;
        RECT 4.400 99.640 146.000 100.960 ;
        RECT 4.400 99.600 145.600 99.640 ;
        RECT 4.000 98.240 145.600 99.600 ;
        RECT 4.000 97.600 146.000 98.240 ;
        RECT 4.400 96.920 146.000 97.600 ;
        RECT 4.400 96.200 145.600 96.920 ;
        RECT 4.000 95.520 145.600 96.200 ;
        RECT 4.000 94.200 146.000 95.520 ;
        RECT 4.400 92.800 145.600 94.200 ;
        RECT 4.000 91.480 146.000 92.800 ;
        RECT 4.000 90.800 145.600 91.480 ;
        RECT 4.400 90.080 145.600 90.800 ;
        RECT 4.400 89.400 146.000 90.080 ;
        RECT 4.000 88.760 146.000 89.400 ;
        RECT 4.000 87.400 145.600 88.760 ;
        RECT 4.400 87.360 145.600 87.400 ;
        RECT 4.400 86.040 146.000 87.360 ;
        RECT 4.400 86.000 145.600 86.040 ;
        RECT 4.000 84.640 145.600 86.000 ;
        RECT 4.000 84.000 146.000 84.640 ;
        RECT 4.400 83.320 146.000 84.000 ;
        RECT 4.400 82.600 145.600 83.320 ;
        RECT 4.000 81.920 145.600 82.600 ;
        RECT 4.000 80.600 146.000 81.920 ;
        RECT 4.400 79.200 145.600 80.600 ;
        RECT 4.000 77.880 146.000 79.200 ;
        RECT 4.000 77.200 145.600 77.880 ;
        RECT 4.400 76.480 145.600 77.200 ;
        RECT 4.400 75.800 146.000 76.480 ;
        RECT 4.000 75.160 146.000 75.800 ;
        RECT 4.000 73.800 145.600 75.160 ;
        RECT 4.400 73.760 145.600 73.800 ;
        RECT 4.400 72.440 146.000 73.760 ;
        RECT 4.400 72.400 145.600 72.440 ;
        RECT 4.000 71.040 145.600 72.400 ;
        RECT 4.000 70.400 146.000 71.040 ;
        RECT 4.400 69.720 146.000 70.400 ;
        RECT 4.400 69.000 145.600 69.720 ;
        RECT 4.000 68.320 145.600 69.000 ;
        RECT 4.000 67.000 146.000 68.320 ;
        RECT 4.400 65.600 145.600 67.000 ;
        RECT 4.000 64.280 146.000 65.600 ;
        RECT 4.000 63.600 145.600 64.280 ;
        RECT 4.400 62.880 145.600 63.600 ;
        RECT 4.400 62.200 146.000 62.880 ;
        RECT 4.000 61.560 146.000 62.200 ;
        RECT 4.000 60.200 145.600 61.560 ;
        RECT 4.400 60.160 145.600 60.200 ;
        RECT 4.400 58.840 146.000 60.160 ;
        RECT 4.400 58.800 145.600 58.840 ;
        RECT 4.000 57.440 145.600 58.800 ;
        RECT 4.000 56.800 146.000 57.440 ;
        RECT 4.400 56.120 146.000 56.800 ;
        RECT 4.400 55.400 145.600 56.120 ;
        RECT 4.000 54.720 145.600 55.400 ;
        RECT 4.000 53.400 146.000 54.720 ;
        RECT 4.400 52.000 145.600 53.400 ;
        RECT 4.000 50.680 146.000 52.000 ;
        RECT 4.000 50.000 145.600 50.680 ;
        RECT 4.400 49.280 145.600 50.000 ;
        RECT 4.400 48.600 146.000 49.280 ;
        RECT 4.000 47.960 146.000 48.600 ;
        RECT 4.000 46.600 145.600 47.960 ;
        RECT 4.400 46.560 145.600 46.600 ;
        RECT 4.400 45.240 146.000 46.560 ;
        RECT 4.400 45.200 145.600 45.240 ;
        RECT 4.000 43.840 145.600 45.200 ;
        RECT 4.000 43.200 146.000 43.840 ;
        RECT 4.400 42.520 146.000 43.200 ;
        RECT 4.400 41.800 145.600 42.520 ;
        RECT 4.000 41.120 145.600 41.800 ;
        RECT 4.000 39.800 146.000 41.120 ;
        RECT 4.400 38.400 145.600 39.800 ;
        RECT 4.000 37.080 146.000 38.400 ;
        RECT 4.000 36.400 145.600 37.080 ;
        RECT 4.400 35.680 145.600 36.400 ;
        RECT 4.400 35.000 146.000 35.680 ;
        RECT 4.000 34.360 146.000 35.000 ;
        RECT 4.000 33.000 145.600 34.360 ;
        RECT 4.400 32.960 145.600 33.000 ;
        RECT 4.400 31.640 146.000 32.960 ;
        RECT 4.400 31.600 145.600 31.640 ;
        RECT 4.000 30.240 145.600 31.600 ;
        RECT 4.000 29.600 146.000 30.240 ;
        RECT 4.400 28.920 146.000 29.600 ;
        RECT 4.400 28.200 145.600 28.920 ;
        RECT 4.000 27.520 145.600 28.200 ;
        RECT 4.000 26.200 146.000 27.520 ;
        RECT 4.400 24.800 145.600 26.200 ;
        RECT 4.000 23.480 146.000 24.800 ;
        RECT 4.000 22.800 145.600 23.480 ;
        RECT 4.400 22.080 145.600 22.800 ;
        RECT 4.400 21.400 146.000 22.080 ;
        RECT 4.000 20.760 146.000 21.400 ;
        RECT 4.000 19.400 145.600 20.760 ;
        RECT 4.400 19.360 145.600 19.400 ;
        RECT 4.400 18.040 146.000 19.360 ;
        RECT 4.400 18.000 145.600 18.040 ;
        RECT 4.000 16.640 145.600 18.000 ;
        RECT 4.000 16.000 146.000 16.640 ;
        RECT 4.400 15.320 146.000 16.000 ;
        RECT 4.400 14.600 145.600 15.320 ;
        RECT 4.000 13.920 145.600 14.600 ;
        RECT 4.000 12.600 146.000 13.920 ;
        RECT 4.400 11.200 146.000 12.600 ;
        RECT 4.000 9.200 146.000 11.200 ;
        RECT 4.400 7.800 146.000 9.200 ;
        RECT 4.000 5.800 146.000 7.800 ;
        RECT 4.400 4.935 146.000 5.800 ;
  END
END tiny_user_project
END LIBRARY

