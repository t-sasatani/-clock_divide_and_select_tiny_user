magic
tech sky130A
magscale 1 2
timestamp 1672324927
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 842 2128 29048 27792
<< metal2 >>
rect 570 29200 626 30000
rect 1674 29200 1730 30000
rect 2778 29200 2834 30000
rect 3882 29200 3938 30000
rect 4986 29200 5042 30000
rect 6090 29200 6146 30000
rect 7194 29200 7250 30000
rect 8298 29200 8354 30000
rect 9402 29200 9458 30000
rect 10506 29200 10562 30000
rect 11610 29200 11666 30000
rect 12714 29200 12770 30000
rect 13818 29200 13874 30000
rect 14922 29200 14978 30000
rect 16026 29200 16082 30000
rect 17130 29200 17186 30000
rect 18234 29200 18290 30000
rect 19338 29200 19394 30000
rect 20442 29200 20498 30000
rect 21546 29200 21602 30000
rect 22650 29200 22706 30000
rect 23754 29200 23810 30000
rect 24858 29200 24914 30000
rect 25962 29200 26018 30000
rect 27066 29200 27122 30000
rect 28170 29200 28226 30000
rect 29274 29200 29330 30000
<< obsm2 >>
rect 682 29144 1618 29322
rect 1786 29144 2722 29322
rect 2890 29144 3826 29322
rect 3994 29144 4930 29322
rect 5098 29144 6034 29322
rect 6202 29144 7138 29322
rect 7306 29144 8242 29322
rect 8410 29144 9346 29322
rect 9514 29144 10450 29322
rect 10618 29144 11554 29322
rect 11722 29144 12658 29322
rect 12826 29144 13762 29322
rect 13930 29144 14866 29322
rect 15034 29144 15970 29322
rect 16138 29144 17074 29322
rect 17242 29144 18178 29322
rect 18346 29144 19282 29322
rect 19450 29144 20386 29322
rect 20554 29144 21490 29322
rect 21658 29144 22594 29322
rect 22762 29144 23698 29322
rect 23866 29144 24802 29322
rect 24970 29144 25906 29322
rect 26074 29144 27010 29322
rect 27178 29144 28114 29322
rect 28282 29144 29042 29322
rect 626 983 29042 29144
<< metal3 >>
rect 0 28840 800 28960
rect 0 28160 800 28280
rect 0 27480 800 27600
rect 0 26800 800 26920
rect 29200 26800 30000 26920
rect 0 26120 800 26240
rect 29200 26256 30000 26376
rect 29200 25712 30000 25832
rect 0 25440 800 25560
rect 29200 25168 30000 25288
rect 0 24760 800 24880
rect 29200 24624 30000 24744
rect 0 24080 800 24200
rect 29200 24080 30000 24200
rect 0 23400 800 23520
rect 29200 23536 30000 23656
rect 29200 22992 30000 23112
rect 0 22720 800 22840
rect 29200 22448 30000 22568
rect 0 22040 800 22160
rect 29200 21904 30000 22024
rect 0 21360 800 21480
rect 29200 21360 30000 21480
rect 0 20680 800 20800
rect 29200 20816 30000 20936
rect 29200 20272 30000 20392
rect 0 20000 800 20120
rect 29200 19728 30000 19848
rect 0 19320 800 19440
rect 29200 19184 30000 19304
rect 0 18640 800 18760
rect 29200 18640 30000 18760
rect 0 17960 800 18080
rect 29200 18096 30000 18216
rect 29200 17552 30000 17672
rect 0 17280 800 17400
rect 29200 17008 30000 17128
rect 0 16600 800 16720
rect 29200 16464 30000 16584
rect 0 15920 800 16040
rect 29200 15920 30000 16040
rect 0 15240 800 15360
rect 29200 15376 30000 15496
rect 29200 14832 30000 14952
rect 0 14560 800 14680
rect 29200 14288 30000 14408
rect 0 13880 800 14000
rect 29200 13744 30000 13864
rect 0 13200 800 13320
rect 29200 13200 30000 13320
rect 0 12520 800 12640
rect 29200 12656 30000 12776
rect 29200 12112 30000 12232
rect 0 11840 800 11960
rect 29200 11568 30000 11688
rect 0 11160 800 11280
rect 29200 11024 30000 11144
rect 0 10480 800 10600
rect 29200 10480 30000 10600
rect 0 9800 800 9920
rect 29200 9936 30000 10056
rect 29200 9392 30000 9512
rect 0 9120 800 9240
rect 29200 8848 30000 8968
rect 0 8440 800 8560
rect 29200 8304 30000 8424
rect 0 7760 800 7880
rect 29200 7760 30000 7880
rect 0 7080 800 7200
rect 29200 7216 30000 7336
rect 29200 6672 30000 6792
rect 0 6400 800 6520
rect 29200 6128 30000 6248
rect 0 5720 800 5840
rect 29200 5584 30000 5704
rect 0 5040 800 5160
rect 29200 5040 30000 5160
rect 0 4360 800 4480
rect 29200 4496 30000 4616
rect 29200 3952 30000 4072
rect 0 3680 800 3800
rect 29200 3408 30000 3528
rect 0 3000 800 3120
rect 29200 2864 30000 2984
rect 0 2320 800 2440
rect 0 1640 800 1760
rect 0 960 800 1080
<< obsm3 >>
rect 880 28080 29200 28253
rect 800 27680 29200 28080
rect 880 27400 29200 27680
rect 800 27000 29200 27400
rect 880 26720 29120 27000
rect 800 26456 29200 26720
rect 800 26320 29120 26456
rect 880 26176 29120 26320
rect 880 26040 29200 26176
rect 800 25912 29200 26040
rect 800 25640 29120 25912
rect 880 25632 29120 25640
rect 880 25368 29200 25632
rect 880 25360 29120 25368
rect 800 25088 29120 25360
rect 800 24960 29200 25088
rect 880 24824 29200 24960
rect 880 24680 29120 24824
rect 800 24544 29120 24680
rect 800 24280 29200 24544
rect 880 24000 29120 24280
rect 800 23736 29200 24000
rect 800 23600 29120 23736
rect 880 23456 29120 23600
rect 880 23320 29200 23456
rect 800 23192 29200 23320
rect 800 22920 29120 23192
rect 880 22912 29120 22920
rect 880 22648 29200 22912
rect 880 22640 29120 22648
rect 800 22368 29120 22640
rect 800 22240 29200 22368
rect 880 22104 29200 22240
rect 880 21960 29120 22104
rect 800 21824 29120 21960
rect 800 21560 29200 21824
rect 880 21280 29120 21560
rect 800 21016 29200 21280
rect 800 20880 29120 21016
rect 880 20736 29120 20880
rect 880 20600 29200 20736
rect 800 20472 29200 20600
rect 800 20200 29120 20472
rect 880 20192 29120 20200
rect 880 19928 29200 20192
rect 880 19920 29120 19928
rect 800 19648 29120 19920
rect 800 19520 29200 19648
rect 880 19384 29200 19520
rect 880 19240 29120 19384
rect 800 19104 29120 19240
rect 800 18840 29200 19104
rect 880 18560 29120 18840
rect 800 18296 29200 18560
rect 800 18160 29120 18296
rect 880 18016 29120 18160
rect 880 17880 29200 18016
rect 800 17752 29200 17880
rect 800 17480 29120 17752
rect 880 17472 29120 17480
rect 880 17208 29200 17472
rect 880 17200 29120 17208
rect 800 16928 29120 17200
rect 800 16800 29200 16928
rect 880 16664 29200 16800
rect 880 16520 29120 16664
rect 800 16384 29120 16520
rect 800 16120 29200 16384
rect 880 15840 29120 16120
rect 800 15576 29200 15840
rect 800 15440 29120 15576
rect 880 15296 29120 15440
rect 880 15160 29200 15296
rect 800 15032 29200 15160
rect 800 14760 29120 15032
rect 880 14752 29120 14760
rect 880 14488 29200 14752
rect 880 14480 29120 14488
rect 800 14208 29120 14480
rect 800 14080 29200 14208
rect 880 13944 29200 14080
rect 880 13800 29120 13944
rect 800 13664 29120 13800
rect 800 13400 29200 13664
rect 880 13120 29120 13400
rect 800 12856 29200 13120
rect 800 12720 29120 12856
rect 880 12576 29120 12720
rect 880 12440 29200 12576
rect 800 12312 29200 12440
rect 800 12040 29120 12312
rect 880 12032 29120 12040
rect 880 11768 29200 12032
rect 880 11760 29120 11768
rect 800 11488 29120 11760
rect 800 11360 29200 11488
rect 880 11224 29200 11360
rect 880 11080 29120 11224
rect 800 10944 29120 11080
rect 800 10680 29200 10944
rect 880 10400 29120 10680
rect 800 10136 29200 10400
rect 800 10000 29120 10136
rect 880 9856 29120 10000
rect 880 9720 29200 9856
rect 800 9592 29200 9720
rect 800 9320 29120 9592
rect 880 9312 29120 9320
rect 880 9048 29200 9312
rect 880 9040 29120 9048
rect 800 8768 29120 9040
rect 800 8640 29200 8768
rect 880 8504 29200 8640
rect 880 8360 29120 8504
rect 800 8224 29120 8360
rect 800 7960 29200 8224
rect 880 7680 29120 7960
rect 800 7416 29200 7680
rect 800 7280 29120 7416
rect 880 7136 29120 7280
rect 880 7000 29200 7136
rect 800 6872 29200 7000
rect 800 6600 29120 6872
rect 880 6592 29120 6600
rect 880 6328 29200 6592
rect 880 6320 29120 6328
rect 800 6048 29120 6320
rect 800 5920 29200 6048
rect 880 5784 29200 5920
rect 880 5640 29120 5784
rect 800 5504 29120 5640
rect 800 5240 29200 5504
rect 880 4960 29120 5240
rect 800 4696 29200 4960
rect 800 4560 29120 4696
rect 880 4416 29120 4560
rect 880 4280 29200 4416
rect 800 4152 29200 4280
rect 800 3880 29120 4152
rect 880 3872 29120 3880
rect 880 3608 29200 3872
rect 880 3600 29120 3608
rect 800 3328 29120 3600
rect 800 3200 29200 3328
rect 880 3064 29200 3200
rect 880 2920 29120 3064
rect 800 2784 29120 2920
rect 800 2520 29200 2784
rect 880 2240 29200 2520
rect 800 1840 29200 2240
rect 880 1560 29200 1840
rect 800 1160 29200 1560
rect 880 987 29200 1160
<< metal4 >>
rect 4417 2128 4737 27792
rect 7890 2128 8210 27792
rect 11363 2128 11683 27792
rect 14836 2128 15156 27792
rect 18309 2128 18629 27792
rect 21782 2128 22102 27792
rect 25255 2128 25575 27792
rect 28728 2128 29048 27792
<< labels >>
rlabel metal3 s 29200 2864 30000 2984 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 29200 19184 30000 19304 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 29200 20816 30000 20936 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 29200 22448 30000 22568 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 29200 24080 30000 24200 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 29200 25712 30000 25832 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 29274 29200 29330 30000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 25962 29200 26018 30000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 22650 29200 22706 30000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 19338 29200 19394 30000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 16026 29200 16082 30000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 29200 4496 30000 4616 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 12714 29200 12770 30000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 9402 29200 9458 30000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 6090 29200 6146 30000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 2778 29200 2834 30000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 29200 6128 30000 6248 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 29200 7760 30000 7880 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 29200 9392 30000 9512 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 29200 11024 30000 11144 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 29200 12656 30000 12776 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 29200 14288 30000 14408 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 29200 15920 30000 16040 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 29200 17552 30000 17672 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 29200 3952 30000 4072 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 29200 20272 30000 20392 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 29200 21904 30000 22024 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 29200 23536 30000 23656 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 29200 25168 30000 25288 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 29200 26800 30000 26920 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 27066 29200 27122 30000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 23754 29200 23810 30000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 20442 29200 20498 30000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 17130 29200 17186 30000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 13818 29200 13874 30000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 29200 5584 30000 5704 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 10506 29200 10562 30000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 7194 29200 7250 30000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 3882 29200 3938 30000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 570 29200 626 30000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 29200 7216 30000 7336 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 960 800 1080 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 29200 8848 30000 8968 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 29200 10480 30000 10600 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 29200 12112 30000 12232 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 29200 13744 30000 13864 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 29200 15376 30000 15496 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 29200 17008 30000 17128 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 29200 18640 30000 18760 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 29200 3408 30000 3528 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 29200 19728 30000 19848 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 29200 21360 30000 21480 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 29200 22992 30000 23112 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 29200 24624 30000 24744 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 29200 26256 30000 26376 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 28170 29200 28226 30000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 24858 29200 24914 30000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 21546 29200 21602 30000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 18234 29200 18290 30000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 14922 29200 14978 30000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 29200 5040 30000 5160 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 11610 29200 11666 30000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 8298 29200 8354 30000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 4986 29200 5042 30000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 1674 29200 1730 30000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 28160 800 28280 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 29200 6672 30000 6792 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 29200 8304 30000 8424 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 29200 9936 30000 10056 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 29200 11568 30000 11688 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 29200 13200 30000 13320 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 29200 14832 30000 14952 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 29200 16464 30000 16584 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 29200 18096 30000 18216 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 4417 2128 4737 27792 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 27792 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 27792 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 27792 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 7890 2128 8210 27792 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 14836 2128 15156 27792 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 21782 2128 22102 27792 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 28728 2128 29048 27792 6 vssd1
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 453344
string GDS_FILE /home/runner/work/clock_divide_and_select_tiny_user/clock_divide_and_select_tiny_user/openlane/tiny_user_project/runs/22_12_29_14_40/results/signoff/tiny_user_project.magic.gds
string GDS_START 23768
<< end >>

